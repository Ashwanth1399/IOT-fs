interface interf ();
  logic clk;
  logic reset;
  logic clear;
  logic [7:0] din;
  logic [7:0] dout;
  logic wr_en;
  logic rd_en;
  logic full;
  logic empty1;

endinterface