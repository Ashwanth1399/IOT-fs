class write_monitor extends uvm_monitor;

  `uvm_component_utils(write_monitor)

  uvm_analysis_port #(fifo_write_sequence_item) item_collected_port_1;

  virtual interf vintf;
  fifo_write_sequence_item fifo_trans;

  function new(string name, uvm_component parent);
    super.new(name, parent);
    fifo_trans = new();
    item_collected_port_1 = new("item_collected_port_1", this);
  endfunction

  function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    fifo_trans = fifo_write_sequence_item::type_id::create("fifo_trans");
    if (!uvm_config_db#(virtual interf)::get(this, "", "vintf", vintf)) begin
      `uvm_error("", "uvm_get_config interface failed\n");
    end
  endfunction

  virtual task run_phase(uvm_phase phase);
    super.run_phase(phase);
    begin
      forever begin
        @(posedge vintf.clk);
        if(vintf.wr_en && !vintf.full) begin
        fifo_trans.wr_en = vintf.wr_en;
        fifo_trans.din   = vintf.din;
        item_collected_port_1.write(fifo_trans);
        `uvm_info("", $sformatf("Monitor: Din is %x\n", vintf.din), UVM_LOW)
        end
      end
    end
  endtask
endclass

